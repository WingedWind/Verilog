module tb;
  // initial begin
  //   $display("Hello from testbench!");
  //   #100;
  //   $display("Bye!");
  //   $finish;
  // end
endmodule